//-----------------------------------------------------------------------------
//  
// MIT License
// Copyright (c) 2022 Advanced Micro Devices, Inc. All rights reserved.
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// SOFTWARE.
//

`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////
// Module Name: xup_and_tb
///////////////////////////////////////////////////////////////

module xup_and_tb(
    );
    
    reg ain, bin;
    reg [2:0] ain_1, bin_1;
    wire y;
    wire [2:0] y_1;
    
    design_1_wrapper DUT(.a(ain), .a_0(ain_1), .b(bin), .b_0(bin_1), .y(y), .y_0(y_1));
    
 
    initial
    begin
      ain = 0; bin= 0; ain_1 = 0; bin_1 = 0;
      #10 ain= 1;
      #10 bin= 1;
	 #10 ain_1 = 3;
	 #10 bin_1 = 1;
      #10 ain= 0; bin= 1;
	 #10 ain_1 = 1; bin_1 = 3;
      #10 ain= 1; bin= 0;
	 #10 ain_1 = 0;
      #10 ain= 1; bin= 1;
      #10 ain= 1; bin= 0;
	#20;
    end

endmodule
